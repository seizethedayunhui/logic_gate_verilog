library verilog;
use verilog.vl_types.all;
entity SnakeTop_tb is
end SnakeTop_tb;
