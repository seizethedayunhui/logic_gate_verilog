library verilog;
use verilog.vl_types.all;
entity tb_Keypad is
end tb_Keypad;
