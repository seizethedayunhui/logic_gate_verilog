library verilog;
use verilog.vl_types.all;
entity tb_StopWatch is
end tb_StopWatch;
