library verilog;
use verilog.vl_types.all;
entity tb_DotMatrixTop is
end tb_DotMatrixTop;
