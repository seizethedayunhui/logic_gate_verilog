library verilog;
use verilog.vl_types.all;
entity tb_logic_test is
end tb_logic_test;
