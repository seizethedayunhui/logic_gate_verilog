library verilog;
use verilog.vl_types.all;
entity tb_UART is
end tb_UART;
