library verilog;
use verilog.vl_types.all;
entity tb_DotMatrix is
end tb_DotMatrix;
