library verilog;
use verilog.vl_types.all;
entity tb_GenEvenParity is
end tb_GenEvenParity;
