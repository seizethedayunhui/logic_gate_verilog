library verilog;
use verilog.vl_types.all;
entity tb_FND is
end tb_FND;
