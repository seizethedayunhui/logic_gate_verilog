library verilog;
use verilog.vl_types.all;
entity tb_SnakeTop is
end tb_SnakeTop;
